library ieee;
use ieee.std_logic_1164.all;

package irig_b_pack is
	constant c_init : std_logic := '1';
	constant c_norm : std_logic := '0';
	
	constant c_frame_size : integer := 10;
end package irig_b_pack;

package body irig_b_pack is

end package body irig_b_pack;
